{\rtf1\ansi\ansicpg936\cocoartf1671\cocoasubrtf400
{\fonttbl\f0\froman\fcharset0 Times-Roman;\f1\fnil\fcharset0 Verdana;}
{\colortbl;\red255\green255\blue255;\red0\green0\blue0;\red255\green255\blue255;}
{\*\expandedcolortbl;;\cssrgb\c0\c0\c0;\cssrgb\c100000\c100000\c100000;}
\paperw11900\paperh16840\margl1440\margr1440\vieww10800\viewh8400\viewkind0
\deftab720
\pard\pardeftab720\sl400\partightenfactor0

\f0\fs28 \cf2 \cb3 \expnd0\expndtw0\kerning0
\
\pard\pardeftab720\sl340\partightenfactor0

\f1 \cf2 module cpu(\cb1 \uc0\u8232 \cb3 \'a0SWB,\cb1 \uc0\u8232 \cb3 \'a0SWA,\cb1 \uc0\u8232 \cb3 \'a0SWC,\cb1 \uc0\u8232 \cb3 \'a0clr,\cb1 \uc0\u8232 \cb3 \'a0C,\cb1 \uc0\u8232 \cb3 \'a0Z,\cb1 \uc0\u8232 \cb3 \'a0IRH,\cb1 \uc0\u8232 \cb3 \'a0T3,\cb1 \uc0\u8232 \cb3 \'a0W1,\cb1 \uc0\u8232 \cb3 \'a0W2,\cb1 \uc0\u8232 \cb3 \'a0W3,\cb1 \uc0\u8232 \cb3 \'a0SELCTL,\cb1 \uc0\u8232 \cb3 \'a0ABUS,\cb1 \uc0\u8232 \cb3 \'a0M,\cb1 \uc0\u8232 \cb3 \'a0S,\cb1 \uc0\u8232 \cb3 \'a0SEL0,\cb1 \uc0\u8232 \cb3 \'a0SEL1,\cb1 \uc0\u8232 \cb3 \'a0SEL2,\cb1 \uc0\u8232 \cb3 \'a0SEL3,\cb1 \uc0\u8232 \cb3 \'a0DRW,\cb1 \uc0\u8232 \cb3 \'a0SBUS,\cb1 \uc0\u8232 \cb3 \'a0LIR,\cb1 \uc0\u8232 \cb3 \'a0MBUS,\cb1 \uc0\u8232 \cb3 \'a0MEMW,\cb1 \uc0\u8232 \cb3 \'a0LAR,\cb1 \uc0\u8232 \cb3 \'a0ARINC,\cb1 \uc0\u8232 \cb3 \'a0LPC,\cb1 \uc0\u8232 \cb3 \'a0PCINC,\cb1 \uc0\u8232 \cb3 \'a0PCADD,\cb1 \uc0\u8232 \cb3 \'a0CIN,\cb1 \uc0\u8232 \cb3 \'a0LONG,\cb1 \uc0\u8232 \cb3 \'a0SHORT,\cb1 \uc0\u8232 \cb3 \'a0CP1,CP2,CP3,\cb1 \uc0\u8232 \cb3 \'a0QD,\cb1 \uc0\u8232 \cb3 \'a0STOP,\cb1 \uc0\u8232 \cb3 \'a0LDC,\cb1 \uc0\u8232 \cb3 \'a0LDZ,\cb1 \uc0\u8232 \cb3 );\cb1 \uc0\u8232 \cb3 input SWB;\cb1 \uc0\u8232 \cb3 input SWA;\cb1 \uc0\u8232 \cb3 input SWC;\cb1 \uc0\u8232 \cb3 input clr;\cb1 \uc0\u8232 \cb3 input C;\cb1 \uc0\u8232 \cb3 input Z;\cb1 \uc0\u8232 \cb3 input [3:0] IRH;\cb1 \uc0\u8232 \cb3 input T3;\cb1 \uc0\u8232 \cb3 input W1;\cb1 \uc0\u8232 \cb3 input W2;\cb1 \uc0\u8232 \cb3 input W3;\cb1 \uc0\u8232 \cb3 input QD;\cb1 \uc0\u8232 \cb3 output SELCTL;\cb1 \uc0\u8232 \cb3 output ABUS;\cb1 \uc0\u8232 \cb3 output M;\cb1 \uc0\u8232 \cb3 output [3:0] S;\cb1 \uc0\u8232 \cb3 output SEL0;\cb1 \uc0\u8232 \cb3 output SEL1;\cb1 \uc0\u8232 \cb3 output SEL2;\cb1 \uc0\u8232 \cb3 output SEL3;\cb1 \uc0\u8232 \cb3 output DRW;\cb1 \uc0\u8232 \cb3 output SBUS;\cb1 \uc0\u8232 \cb3 output LIR;\cb1 \uc0\u8232 \cb3 output MBUS;\cb1 \uc0\u8232 \cb3 output MEMW;\cb1 \uc0\u8232 \cb3 output LAR;\cb1 \uc0\u8232 \cb3 output ARINC;\cb1 \uc0\u8232 \cb3 output LPC;\cb1 \uc0\u8232 \cb3 output PCINC;\cb1 \uc0\u8232 \cb3 output PCADD;\cb1 \uc0\u8232 \cb3 output CIN;\cb1 \uc0\u8232 \cb3 output LONG;\cb1 \uc0\u8232 \cb3 output SHORT;\cb1 \uc0\u8232 \cb3 output STOP;\cb1 \uc0\u8232 \cb3 output LDC;\cb1 \uc0\u8232 \cb3 output LDZ;\cb1 \uc0\u8232 \cb3 output CP1,CP2,CP3;\cb1 \uc0\u8232 \cb3 reg SELCTL;\cb1 \uc0\u8232 \cb3 reg ABUS;\cb1 \uc0\u8232 \cb3 reg M;\cb1 \uc0\u8232 \cb3 reg [3:0] S;\cb1 \uc0\u8232 \cb3 reg SEL0;\cb1 \uc0\u8232 \cb3 reg SEL1;\cb1 \uc0\u8232 \cb3 reg SEL2;\cb1 \uc0\u8232 \cb3 reg SEL3;\cb1 \uc0\u8232 \cb3 reg DRW;\cb1 \uc0\u8232 \cb3 reg SBUS;\cb1 \uc0\u8232 \cb3 reg LIR;\cb1 \uc0\u8232 \cb3 reg MBUS;\cb1 \uc0\u8232 \cb3 reg MEMW;\cb1 \uc0\u8232 \cb3 reg LAR;\cb1 \uc0\u8232 \cb3 reg ARINC;\cb1 \uc0\u8232 \cb3 reg LPC;\cb1 \uc0\u8232 \cb3 reg PCINC;\cb1 \uc0\u8232 \cb3 reg PCADD;\cb1 \uc0\u8232 \cb3 reg CIN;\cb1 \uc0\u8232 \cb3 reg LONG;\cb1 \uc0\u8232 \cb3 reg SHORT;\cb1 \uc0\u8232 \cb3 reg LDC;\cb1 \uc0\u8232 \cb3 reg LDZ;\cb1 \uc0\u8232 \cb3 wire[2:0] SWCBA;\cb1 \uc0\u8232 \cb3 wire ST0;\cb1 \uc0\u8232 \cb3 wire ST1;\cb1 \uc0\u8232 \cb3 reg ST0_reg;\cb1 \uc0\u8232 \cb3 reg ST1_reg;\cb1 \uc0\u8232 \cb3 reg SST0;\cb1 \uc0\u8232 \cb3 reg SST1;\cb1 \uc0\u8232 \cb3 wire STOP;\cb1 \uc0\u8232 \cb3 reg STOP_reg_reg_reg;\cb1 \uc0\u8232 \cb3 reg STOP_reg_reg;\cb1 \uc0\u8232 \cb3 reg STOP_reg;\cb1 \uc0\u8232 \cb3 parameter\cb1 \uc0\u8232 \cb3 NOP=4'B0000,\cb1 \uc0\u8232 \cb3 ADD=4'b0001,\cb1 \uc0\u8232 \cb3 SUB=4'B0010,\cb1 \uc0\u8232 \cb3 AND=4'B0011,\cb1 \uc0\u8232 \cb3 INC=4'B0100,\cb1 \uc0\u8232 \cb3 LD=4'B0101,\cb1 \uc0\u8232 \cb3 ST=4'B0110,\cb1 \uc0\u8232 \cb3 JC=4'B0111,\cb1 \uc0\u8232 \cb3 JZ=4'B1000,\cb1 \uc0\u8232 \cb3 JMP=4'B1001,\cb1 \uc0\u8232 \cb3 OUT=4'B1010,\cb1 \uc0\u8232 \cb3 STP=4'B1110,\cb1 \uc0\u8232 \cb3 OR=4'B1011,\cb1 \uc0\u8232 \cb3 XAND=4'B1100,\cb1 \uc0\u8232 \cb3 LSHIFT=4'B1101;\cb1 \uc0\u8232 \cb3 assign STOP=(SWCBA?(STOP_reg_reg|STOP_reg|STOP_reg_reg_reg):0);\cb1 \uc0\u8232 \cb3 assign CP1=1'b1;\cb1 \uc0\u8232 \cb3 assign CP2=1'b1;\cb1 \uc0\u8232 \cb3 assign CP3=QD;\cb1 \uc0\u8232 \cb3 assign SWCBA[2:0]=\{SWC,SWB,SWA\};\cb1 \uc0\u8232 \cb3 assign ST0=ST0_reg;\cb1 \uc0\u8232 \cb3 assign ST1=ST1_reg;\cb1 \uc0\u8232 \cb3 always @(negedge clr or negedge T3)\cb1 \uc0\u8232 \cb3 begin\cb1 \uc0\u8232 \cb3 \'a0if(clr==0)\cb1 \uc0\u8232 \cb3 \'a0begin\cb1 \uc0\u8232 \cb3 \'a0 ST0_reg<=0;\cb1 \uc0\u8232 \cb3 \'a0 STOP_reg_reg<=1;\cb1 \uc0\u8232 \cb3 \'a0end\cb1 \uc0\u8232 \cb3 \'a0else\cb1 \uc0\u8232 \cb3 \'a0begin\cb1 \uc0\u8232 \cb3 \'a0 if(SST0==1'b1) ST0_reg<=1'b1;\cb1 \uc0\u8232 \cb3 \'a0end\cb1 \uc0\u8232 \cb3 end
\f0 \

\f1 always @(negedge clr or negedge T3)\cb1 \uc0\u8232 \cb3 begin\cb1 \uc0\u8232 \cb3 \'a0if(clr==0)\cb1 \uc0\u8232 \cb3 \'a0begin\cb1 \uc0\u8232 \cb3 \'a0 ST1_reg<=0;\cb1 \uc0\u8232 \cb3 \'a0 STOP_reg_reg_reg<=1;\cb1 \uc0\u8232 \cb3 \'a0end\cb1 \uc0\u8232 \cb3 \'a0else\cb1 \uc0\u8232 \cb3 \'a0begin\cb1 \uc0\u8232 \cb3 \'a0 if((SST1==1'b1)&(ST1_reg==1'b0)) ST1_reg<=1'b1;\cb1 \uc0\u8232 \cb3 \'a0 else if((SST1==1'b1)&(ST1_reg==1'b1)) ST1_reg<=1'b0;\cb1 \uc0\u8232 \cb3 \'a0end\cb1 \uc0\u8232 \cb3 end
\f0 \

\f1 always @ (W1 or W2 or W3 or ST0 or C or Z or SWCBA or IRH)\cb1 \uc0\u8232 \cb3 begin\cb1 \uc0\u8232 \cb3 \'a0SELCTL <=0;\cb1 \uc0\u8232 \cb3 \'a0ABUS\'a0 <=0;\cb1 \uc0\u8232 \cb3 \'a0M \'a0 <=0;\cb1 \uc0\u8232 \cb3 \'a0S \'a0 <=4'b0000;\cb1 \uc0\u8232 \cb3 \'a0SEL0\'a0 <=0;\cb1 \uc0\u8232 \cb3 \'a0SEL1\'a0 <=0;\cb1 \uc0\u8232 \cb3 \'a0SEL2\'a0 <=0;\cb1 \uc0\u8232 \cb3 \'a0SEL3\'a0 <=0;\cb1 \uc0\u8232 \cb3 \'a0DRW\'a0\'a0\'a0 \'a0 <=0;\cb1 \uc0\u8232 \cb3 \'a0SBUS\'a0 <=0;\cb1 \uc0\u8232 \cb3 \'a0LIR\'a0\'a0\'a0 \'a0 <=0;\cb1 \uc0\u8232 \cb3 \'a0MBUS\'a0 <=0;\cb1 \uc0\u8232 \cb3 \'a0MEMW\'a0 <=0;\cb1 \uc0\u8232 \cb3 \'a0LAR\'a0\'a0\'a0 \'a0 <=0;\cb1 \uc0\u8232 \cb3 \'a0ARINC\'a0 <=0;\cb1 \uc0\u8232 \cb3 \'a0LPC\'a0\'a0\'a0 \'a0 <=0;\cb1 \uc0\u8232 \cb3 \'a0PCINC\'a0 <=0;\cb1 \uc0\u8232 \cb3 \'a0CIN\'a0\'a0\'a0 \'a0 <=0;\cb1 \uc0\u8232 \cb3 \'a0LONG\'a0 <=0;\cb1 \uc0\u8232 \cb3 \'a0SHORT\'a0 <=0;\cb1 \uc0\u8232 \cb3 \'a0LDZ\'a0\'a0\'a0 \'a0 <=0;\cb1 \uc0\u8232 \cb3 \'a0LDC\'a0\'a0\'a0 \'a0 <=0;\cb1 \uc0\u8232 \cb3 \'a0PCADD\'a0 <=0;\cb1 \uc0\u8232 \cb3 \'a0STOP_reg <=1;\cb1 \uc0\u8232 \cb3 \'a0SST0\'a0 <=0;\cb1 \uc0\u8232 \cb3 \'a0\cb1 \uc0\u8232 \cb3 \'a0case(SWCBA)\cb1 \uc0\u8232 \cb3 \'a0 3'b000:\cb1 \uc0\u8232 \cb3 \'a0 begin\cb1 \uc0\u8232 \cb3 \'a0\'a0 if(ST0==0)\cb1 \uc0\u8232 \cb3 \'a0 \'a0 begin\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 SBUS<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 LPC<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 SHORT<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 SST0<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 STOP_reg<=0;\cb1 \uc0\u8232 \cb3 \'a0 \'a0 end\cb1 \uc0\u8232 \cb3 \'a0\'a0 else if(ST0==1)\cb1 \uc0\u8232 \cb3 \'a0 \'a0 begin\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 case(IRH)\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0 \'a0 NOP:\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 begin\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LIR<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 PCINC<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 SHORT<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 end\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0 \'a0 ADD:\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 begin\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 CIN<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 ABUS<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 DRW<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LDZ<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LDC<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 S<=4'b1001;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0\'a0\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LIR<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 PCINC<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 SHORT<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 end\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0 \'a0 SUB:\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 begin\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 ABUS<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 DRW<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LDZ<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LDC<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 S<=4'b0110;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0\'a0\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LIR<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 PCINC<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 SHORT<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 end\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0 \'a0 AND:\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 begin\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 M<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 ABUS<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 DRW<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LDZ<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 S<=4'B1011;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0\'a0\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LIR<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 PCINC<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 SHORT<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 end\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0 \'a0 INC:\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 begin\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 ABUS<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 DRW<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LDZ<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LDC<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 S<=4'B0000;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0\'a0\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LIR<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 PCINC<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 SHORT<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 end\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0 \'a0 LD:\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 begin\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 M<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 ABUS<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LAR<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 S<=4'B1010;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 MBUS<=W2;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 DRW<=W2;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0\'a0\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LIR<=W2;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 PCINC<=W2;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 end\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0 \'a0 ST:\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 begin\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 M<=W1|W2;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 ABUS<=W2|W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LAR<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 S[3]<=1'B1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 S[1]<=1'B1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 S[2]<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 S[0]<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 MEMW<=W2;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0\'a0\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LIR<=W2;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 PCINC<=W2;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 end\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0 \'a0 JC:\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 begin\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 PCADD<=C&W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0\'a0\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LIR<=(W1&(~C))|(W2&C);\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 PCINC<=(W1&(~C))|(W2&C);\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 SHORT<=W1&(~C);\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 end\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0 \'a0 JZ:\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 begin\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 PCADD<=Z&W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0\'a0\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LIR<=(W1&(~Z))|(W2&Z);\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 PCINC<=(W1&(~Z))|(W2&Z);\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 SHORT<=W1&(~Z);\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 end\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0 \'a0 JMP:\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 begin\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 M<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 S<=4'b1111;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 ABUS<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LPC<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0\'a0\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LIR<=W2;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 PCINC<=W2;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 end\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0 \'a0 STP:\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 begin\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 STOP_reg<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 end\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0 \'a0 OUT:\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 begin\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 M<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 S<=4'b1010;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 ABUS<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0\'a0\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LIR<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 PCINC<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 SHORT<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 end\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0 \'a0 OR:\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 begin\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 M<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 ABUS<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 DRW<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LDZ<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 S<=4'b1110;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0\'a0\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LIR<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 PCINC<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 SHORT<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 end\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0 \'a0 XAND:\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 begin\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 M<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 ABUS<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 DRW<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LDZ<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 S<=4'b0100;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0\'a0\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LIR<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 PCINC<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 SHORT<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 end\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0 \'a0 LSHIFT:\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 begin\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 CIN<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 ABUS<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 DRW<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LDZ<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LDC<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 S<=4'b1100;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0\'a0\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 LIR<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 PCINC<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0\'a0 \'a0 SHORT<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 end\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0 \'a0 default:\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 begin\cb1 \uc0\u8232 \cb3 \'a0 LIR<=W1;\cb1 \uc0\u8232 \cb3 \'a0 PCINC<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0\'a0\'a0 \'a0 end\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 endcase\cb1 \uc0\u8232 \cb3 \'a0 \'a0 end\cb1 \uc0\u8232 \cb3 \'a0\'a0 end\cb1 \uc0\u8232 \cb3 \'a0\cb1 \uc0\u8232 \cb3 \'a0\'a0 3'b001:\cb1 \uc0\u8232 \cb3 \'a0 \'a0 begin\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 SELCTL<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 SHORT<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 SBUS<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 STOP_reg<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 SST0<=W1;\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 LAR<=W1&(~ST0);\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 ARINC<=W1&ST0;\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 MEMW<=W1&ST0;\cb1 \uc0\u8232 \cb3 \'a0 \'a0 end\cb1 \uc0\u8232 \cb3 \'a0\cb1 \uc0\u8232 \cb3 \'a0\'a0 3'b011:\cb1 \uc0\u8232 \cb3 \'a0 \'a0 begin\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 SELCTL<=1'b1;\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 SEL0<=W1|W2;\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 STOP_reg<=W1|W2;\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 SEL3<=W2;\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 SEL1<=W2;\cb1 \uc0\u8232 \cb3 \'a0 \'a0 end\cb1 \uc0\u8232 \cb3 \'a0\cb1 \uc0\u8232 \cb3 \'a0\'a0 3'b100:\cb1 \uc0\u8232 \cb3 \'a0 \'a0 begin\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 SELCTL<=1'b1;\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 SST1<=W2;\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 SBUS<=W1|W2;\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 STOP_reg<=W1|W2;\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 DRW<=W1|W2;\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 SEL3<=(ST1&W1)|(ST1&W2);\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 SEL2<=W2;\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 SEL1<=((~ST1)&W1)|(ST1&W2);\cb1 \uc0\u8232 \cb3 \'a0\'a0 \'a0 SEL0<=W1;\cb1 \uc0\u8232 \cb3 \'a0 \'a0 end\cb1 \uc0\u8232 \cb3 \'a0\cb1 \uc0\u8232 \cb3 \'a03'b010:\cb1 \uc0\u8232 \cb3 \'a0 begin\cb1 \uc0\u8232 \cb3 \'a0 SBUS<=(~ST0)&W1;\cb1 \uc0\u8232 \cb3 \'a0 LAR<=(~ST0)&W1;\cb1 \uc0\u8232 \cb3 \'a0 STOP_reg<=W1;\cb1 \uc0\u8232 \cb3 \'a0 SST0<=(~ST0)&W1;\cb1 \uc0\u8232 \cb3 \'a0 SHORT<=W1;\cb1 \uc0\u8232 \cb3 \'a0 SELCTL<=W1;\cb1 \uc0\u8232 \cb3 \'a0 MBUS<=ST0&W1;\cb1 \uc0\u8232 \cb3 \'a0 ARINC<=ST0&W1;\cb1 \uc0\u8232 \cb3 \'a0end\cb1 \uc0\u8232 \cb3 \'a0\'a0\cb1 \uc0\u8232 \cb3 \'a0\'a0 default:\cb1 \uc0\u8232 \cb3 \'a0 \'a0 begin\cb1 \uc0\u8232 \cb3 \'a0 \'a0 end\cb1 \uc0\u8232 \cb3 \'a0endcase\cb1 \uc0\u8232 \cb3 end\cb1 \uc0\u8232 \cb3 endmodule
\f0 \
}