{\rtf1\ansi\ansicpg936\cocoartf1671\cocoasubrtf400
{\fonttbl\f0\fnil\fcharset0 Verdana;\f1\froman\fcharset0 Times-Roman;}
{\colortbl;\red255\green255\blue255;\red0\green0\blue0;\red255\green255\blue255;}
{\*\expandedcolortbl;;\cssrgb\c0\c0\c0;\cssrgb\c100000\c100000\c100000;}
\paperw11900\paperh16840\margl1440\margr1440\vieww10800\viewh8400\viewkind0
\deftab720
\pard\pardeftab720\sl340\sa0\partightenfactor0

\f0\fs28 \cf2 \cb3 \expnd0\expndtw0\kerning0
\outl0\strokewidth0 \strokec2 module CPU(
\f1 \

\f0 \'a0SWB,
\f1 \

\f0 \'a0SWA,
\f1 \

\f0 \'a0SWC,
\f1 \

\f0 \'a0clr,
\f1 \

\f0 \'a0C,
\f1 \

\f0 \'a0Z,
\f1 \

\f0 \'a0IRH,
\f1 \

\f0 \'a0T3,
\f1 \

\f0 \'a0W1,
\f1 \

\f0 \'a0W2,
\f1 \

\f0 \'a0W3,
\f1 \

\f0 \'a0SELCTL,
\f1 \

\f0 \'a0ABUS,
\f1 \

\f0 \'a0M,
\f1 \

\f0 \'a0S,
\f1 \

\f0 \'a0SEL0,
\f1 \

\f0 \'a0SEL1,
\f1 \

\f0 \'a0SEL2,
\f1 \

\f0 \'a0SEL3,
\f1 \

\f0 \'a0DRW,
\f1 \

\f0 \'a0SBUS,
\f1 \

\f0 \'a0LIR,
\f1 \

\f0 \'a0MBUS,
\f1 \

\f0 \'a0MEMW,
\f1 \

\f0 \'a0LAR,
\f1 \

\f0 \'a0ARINC,
\f1 \

\f0 \'a0LPC,
\f1 \

\f0 \'a0PCINC,
\f1 \

\f0 \'a0PCADD,
\f1 \

\f0 \'a0CIN,
\f1 \

\f0 \'a0LONG,
\f1 \

\f0 \'a0SHORT,
\f1 \

\f0 \'a0CP1,CP2,CP3,
\f1 \

\f0 \'a0QD,
\f1 \

\f0 \'a0STOP,
\f1 \

\f0 \'a0LDC,
\f1 \

\f0 \'a0LDZ,
\f1 \

\f0 );
\f1 \

\f0 input SWB;
\f1 \

\f0 input SWA;
\f1 \

\f0 input SWC;
\f1 \

\f0 input clr;
\f1 \

\f0 input C;
\f1 \

\f0 input Z;
\f1 \

\f0 input [3:0] IRH;
\f1 \

\f0 input T3;
\f1 \

\f0 input W1;
\f1 \

\f0 input W2;
\f1 \

\f0 input W3;
\f1 \

\f0 input QD;
\f1 \

\f0 output SELCTL;
\f1 \

\f0 output ABUS;
\f1 \

\f0 output M;
\f1 \

\f0 output [3:0] S;
\f1 \

\f0 output SEL0;
\f1 \

\f0 output SEL1;
\f1 \

\f0 output SEL2;
\f1 \

\f0 output SEL3;
\f1 \

\f0 output DRW;
\f1 \

\f0 output SBUS;
\f1 \

\f0 output LIR;
\f1 \

\f0 output MBUS;
\f1 \

\f0 output MEMW;
\f1 \

\f0 output LAR;
\f1 \

\f0 output ARINC;
\f1 \

\f0 output LPC;
\f1 \

\f0 output PCINC;
\f1 \

\f0 output PCADD;
\f1 \

\f0 output CIN;
\f1 \

\f0 output LONG;
\f1 \

\f0 output SHORT;
\f1 \

\f0 output STOP;
\f1 \

\f0 output LDC;
\f1 \

\f0 output LDZ;
\f1 \

\f0 output CP1,CP2,CP3;
\f1 \

\f0 reg SELCTL;
\f1 \

\f0 reg ABUS;
\f1 \

\f0 reg M;
\f1 \

\f0 reg [3:0] S;
\f1 \

\f0 reg SEL0;
\f1 \

\f0 reg SEL1;
\f1 \

\f0 reg SEL2;
\f1 \

\f0 reg SEL3;
\f1 \

\f0 reg DRW;
\f1 \

\f0 reg SBUS;
\f1 \

\f0 reg LIR;
\f1 \

\f0 reg MBUS;
\f1 \

\f0 reg MEMW;
\f1 \

\f0 reg LAR;
\f1 \

\f0 reg ARINC;
\f1 \

\f0 reg LPC;
\f1 \

\f0 reg PCINC;
\f1 \

\f0 reg PCADD;
\f1 \

\f0 reg CIN;
\f1 \

\f0 reg LONG;
\f1 \

\f0 reg SHORT;
\f1 \

\f0 reg LDC;
\f1 \

\f0 reg LDZ;
\f1 \

\f0 wire[2:0] SWCBA;
\f1 \

\f0 wire ST0;
\f1 \

\f0 wire ST1;
\f1 \

\f0 reg ST0_reg;
\f1 \

\f0 reg ST1_reg;
\f1 \

\f0 reg SST0;
\f1 \

\f0 reg SST1;
\f1 \

\f0 wire STOP;
\f1 \

\f0 reg STOP_reg_reg;
\f1 \

\f0 reg STOP_reg_reg_reg;
\f1 \

\f0 reg STOP_reg;
\f1 \

\f0 parameter 
\f1 \

\f0 ADD=4'b0001,
\f1 \

\f0 SUB=4'B0010,
\f1 \

\f0 AND=4'B0011,
\f1 \

\f0 INC=4'B0100,
\f1 \

\f0 LD=4'B0101,
\f1 \

\f0 ST=4'B0110,
\f1 \

\f0 JC=4'B0111,
\f1 \

\f0 JZ=4'B1000,
\f1 \

\f0 JMP=4'B1001,
\f1 \

\f0 OUT=4'B1010,
\f1 \

\f0 STP=4'B1110,
\f1 \

\f0 OR=4'B1011,
\f1 \

\f0 XAND=4'B1100,
\f1 \

\f0 LSHIFT=4'B1101;
\f1 \

\f0 assign STOP=(SWCBA?(STOP_reg_reg|STOP_reg|STOP_reg_reg_reg):0);
\f1 \

\f0 assign CP1=1'b1;
\f1 \

\f0 assign CP2=1'b1;
\f1 \

\f0 assign CP3=QD;
\f1 \

\f0 assign SWCBA[2:0]=\{SWC,SWB,SWA\};
\f1 \

\f0 assign ST0=ST0_reg;
\f1 \

\f0 assign ST1=ST1_reg;
\f1 \

\f0 always @(negedge clr or negedge T3)
\f1 \

\f0 begin
\f1 \

\f0 \'a0if(clr==0)
\f1 \

\f0 \'a0begin
\f1 \

\f0 \'a0 ST0_reg<=0;
\f1 \

\f0 \'a0 STOP_reg_reg<=1;
\f1 \

\f0 \'a0end
\f1 \

\f0 \'a0else
\f1 \

\f0 \'a0begin
\f1 \

\f0 \'a0 if(SST0==1'b1) ST0_reg<=1'b1;
\f1 \

\f0 \'a0end
\f1 \

\f0 end
\f1 \

\f0 always @(negedge clr or negedge T3)
\f1 \

\f0 begin
\f1 \

\f0 \'a0if(clr==0)
\f1 \

\f0 \'a0begin
\f1 \

\f0 \'a0 ST1_reg<=0;
\f1 \

\f0 \'a0 STOP_reg_reg_reg<=1;
\f1 \

\f0 \'a0end
\f1 \

\f0 \'a0else
\f1 \

\f0 \'a0begin
\f1 \

\f0 \'a0 if((SST1==1'b1)&(ST1_reg==1'b0)) ST1_reg<=1'b1;
\f1 \

\f0 \'a0 else if((SST1==1'b1)&(ST1_reg==1'b1)) ST1_reg<=1'b0;
\f1 \

\f0 \'a0end
\f1 \

\f0 end
\f1 \

\f0 always @ (W1 or W2 or W3 or ST0 or C or Z or SWCBA or IRH)
\f1 \

\f0 begin
\f1 \

\f0 \'a0SELCTL <=0;
\f1 \

\f0 \'a0ABUS\'a0 <=0;
\f1 \

\f0 \'a0M\'a0 \'a0<=0;
\f1 \

\f0 \'a0S\'a0 \'a0<=4'b0000;
\f1 \

\f0 \'a0SEL0\'a0 <=0;
\f1 \

\f0 \'a0SEL1\'a0 <=0;
\f1 \

\f0 \'a0SEL2\'a0 <=0;
\f1 \

\f0 \'a0SEL3\'a0 <=0;
\f1 \

\f0 \'a0DRW\'a0 <=0;
\f1 \

\f0 \'a0SBUS\'a0 <=0;
\f1 \

\f0 \'a0LIR\'a0 <=0;
\f1 \

\f0 \'a0MBUS\'a0 <=0;
\f1 \

\f0 \'a0MEMW\'a0 <=0;
\f1 \

\f0 \'a0LAR\'a0 <=0;
\f1 \

\f0 \'a0ARINC\'a0 <=0;
\f1 \

\f0 \'a0LPC\'a0 <=0;
\f1 \

\f0 \'a0PCINC\'a0 <=0;
\f1 \

\f0 \'a0CIN\'a0 <=0;
\f1 \

\f0 \'a0LONG\'a0 <=0;
\f1 \

\f0 \'a0SHORT\'a0 <=0;
\f1 \

\f0 \'a0LDZ\'a0 <=0;
\f1 \

\f0 \'a0LDC\'a0 <=0;
\f1 \

\f0 \'a0PCADD\'a0 <=0;
\f1 \

\f0 \'a0STOP_reg <=1;
\f1 \

\f0 \'a0SST0\'a0 <=0;
\f1 \

\f0 \'a0SST1\'a0 <=0;
\f1 \

\f0 \'a0
\f1 \

\f0 \'a0case(SWCBA)
\f1 \

\f0 \'a0 3'b000:
\f1 \

\f0 \'a0 begin
\f1 \

\f0 \'a0 \'a0if(ST0==0)
\f1 \

\f0 \'a0 \'a0 begin
\f1 \

\f0 \'a0 \'a0 \'a0SBUS<=W1;
\f1 \

\f0 \'a0 \'a0 \'a0LPC<=W1;
\f1 \

\f0 \'a0 \'a0 \'a0SHORT<=W1;
\f1 \

\f0 \'a0 \'a0 \'a0SST0<=W1;
\f1 \

\f0 \'a0 \'a0 \'a0STOP_reg<=0;
\f1 \

\f0 \'a0 \'a0 end
\f1 \

\f0 \'a0 \'a0else if(ST0==1)
\f1 \

\f0 \'a0 \'a0 begin
\f1 \

\f0 \'a0 \'a0 \'a0LIR<=W1;
\f1 \

\f0 \'a0 \'a0 \'a0PCINC<=W1;
\f1 \

\f0 \'a0 \'a0 \'a0case(IRH)
\f1 \

\f0 \'a0 \'a0 \'a0 ADD:
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0begin
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 CIN<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 ABUS<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 DRW<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 LDZ<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 LDC<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 S<=4'b1001;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0end
\f1 \

\f0 \'a0 \'a0 \'a0 SUB:
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0begin
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 ABUS<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 DRW<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 LDZ<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 LDC<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 S<=4'b0110;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0end
\f1 \

\f0 \'a0 \'a0 \'a0 AND:
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0begin
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 M<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 ABUS<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 DRW<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 LDZ<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 S<=4'B1011;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0end
\f1 \

\f0 \'a0 \'a0 \'a0 INC:
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0begin
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 ABUS<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 DRW<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 LDZ<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 LDC<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 S<=4'B0000;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0end
\f1 \

\f0 \'a0 \'a0 \'a0 LD:
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0begin
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 M<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 ABUS<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 LAR<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 LONG<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 S<=4'B1010;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 MBUS<=W3;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 DRW<=W3;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0end
\f1 \

\f0 \'a0 \'a0 \'a0 ST:
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0begin
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 M<=W2|W3;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 ABUS<=W2|W3;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 LAR<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 LONG<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 S[3]<=1'B1;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 S[1]<=1'B1;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 S[2]<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 S[0]<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 MEMW<=W3;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0end
\f1 \

\f0 \'a0 \'a0 \'a0 JC:
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0begin
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 PCADD<=C&W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0end
\f1 \

\f0 \'a0 \'a0 \'a0 JZ:
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0begin
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 PCADD<=Z&W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0end
\f1 \

\f0 \'a0 \'a0 \'a0 JMP:
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0begin
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 M<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 S<=4'b1111;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 ABUS<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 LPC<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0end
\f1 \

\f0 \'a0 \'a0 \'a0 STP:
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0begin
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 STOP_reg<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0end
\f1 \

\f0 \'a0 \'a0 \'a0 OUT:
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0begin
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 M<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 S<=4'b1010;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 ABUS<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0end
\f1 \

\f0 \'a0 \'a0 \'a0 OR:
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0begin
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 M<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 ABUS<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 DRW<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 LDZ<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 S<=4'B1110;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0end
\f1 \

\f0 \'a0 \'a0 \'a0 XAND:
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0begin
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 M<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 ABUS<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 DRW<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 LDZ<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 S<=4'B0100;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0end
\f1 \

\f0 \'a0 \'a0 \'a0 LSHIFT:
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0begin
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 CIN<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 ABUS<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 DRW<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 LDZ<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 LDC<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0 S<=4'b1100;
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0end
\f1 \

\f0 \'a0 \'a0 \'a0 default:
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0begin
\f1 \

\f0 \'a0 \'a0 \'a0 \'a0end
\f1 \

\f0 \'a0 \'a0 \'a0endcase
\f1 \

\f0 \'a0 \'a0 end
\f1 \

\f0 \'a0 \'a0end
\f1 \

\f0 \'a0
\f1 \

\f0 \'a0 \'a03'b001:
\f1 \

\f0 \'a0 \'a0 begin
\f1 \

\f0 \'a0 \'a0 \'a0SELCTL<=W1;
\f1 \

\f0 \'a0 \'a0 \'a0SHORT<=W1;
\f1 \

\f0 \'a0 \'a0 \'a0SBUS<=W1;
\f1 \

\f0 \'a0 \'a0 \'a0STOP_reg<=W1;
\f1 \

\f0 \'a0 \'a0 \'a0SST0<=W1;
\f1 \

\f0 \'a0 \'a0 \'a0LAR<=W1&(~ST0);
\f1 \

\f0 \'a0 \'a0 \'a0ARINC<=W1&ST0;
\f1 \

\f0 \'a0 \'a0 \'a0MEMW<=W1&ST0;
\f1 \

\f0 \'a0 \'a0 end
\f1 \

\f0 \'a0
\f1 \

\f0 \'a0 \'a03'b011:
\f1 \

\f0 \'a0 \'a0 begin
\f1 \

\f0 \'a0 \'a0 \'a0SELCTL<=1'b1;
\f1 \

\f0 \'a0 \'a0 \'a0SEL0<=W1|W2;
\f1 \

\f0 \'a0 \'a0 \'a0STOP_reg<=W1|W2;
\f1 \

\f0 \'a0 \'a0 \'a0SEL3<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0SEL1<=W2;
\f1 \

\f0 \'a0 \'a0 end
\f1 \

\f0 \'a0
\f1 \

\f0 \'a0 \'a03'b100:
\f1 \

\f0 \'a0 \'a0 begin
\f1 \

\f0 \'a0 \'a0 \'a0SELCTL<=1'b1;
\f1 \

\f0 \'a0 \'a0 \'a0SST1<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0SBUS<=W1|W2;
\f1 \

\f0 \'a0 \'a0 \'a0STOP_reg<=W1|W2;
\f1 \

\f0 \'a0 \'a0 \'a0DRW<=W1|W2;
\f1 \

\f0 \'a0 \'a0 \'a0if(ST1==0)
\f1 \

\f0 \'a0 \'a0 \'a0begin
\f1 \

\f0 \'a0 \'a0 \'a0 SEL1<=W1;
\f1 \

\f0 \'a0 \'a0 \'a0end
\f1 \

\f0 \'a0 \'a0 \'a0else
\f1 \

\f0 \'a0 \'a0 \'a0begin
\f1 \

\f0 \'a0 \'a0 \'a0 SEL3<=W1|W2;
\f1 \

\f0 \'a0 \'a0 \'a0 SEL1<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0end
\f1 \

\f0 \'a0 \'a0 \'a0SEL2<=W2;
\f1 \

\f0 \'a0 \'a0 \'a0SEL0<=W1;
\f1 \

\f0 \'a0 \'a0 end
\f1 \

\f0 \'a0
\f1 \

\f0 \'a0 \'a03'b010:
\f1 \

\f0 \'a0 \'a0 begin
\f1 \

\f0 \'a0 \'a0 \'a0SUBS<=(~ST0)&W1;
\f1 \

\f0 \'a0 \'a0 \'a0LAR<=(~ST0)&W1;
\f1 \

\f0 \'a0 \'a0 \'a0STOP_reg<=W1;
\f1 \

\f0 \'a0 \'a0 \'a0SST0<=(~ST0)&W1;
\f1 \

\f0 \'a0 \'a0 \'a0SHORT<=W1;
\f1 \

\f0 \'a0 \'a0 \'a0SELCTL<=W1;
\f1 \

\f0 \'a0 \'a0 \'a0MUBS<=ST0&W1;
\f1 \

\f0 \'a0 \'a0 \'a0ARINC<=ST0&W1;
\f1 \

\f0 \'a0 \'a0 end
\f1 \

\f0 \'a0
\f1 \

\f0 \'a0 \'a0default:
\f1 \

\f0 \'a0 \'a0 begin
\f1 \

\f0 \'a0 \'a0 end
\f1 \

\f0 \'a0endcase
\f1 \

\f0 end
\f1 \

\f0 endmodule
\f1 \

\f0 \'a0
\f1 \

\f0 \'a0
\f1 \

\f0 \'a0
\f1 \

\f0 \'a0
\f1 \

\f0 \'a0
\f1 \

\f0 \'a0
\f1 \

\f0 \'a0
\f1 \

\f0 \'a0
\f1 \

\f0 \'a0
\f1 \

\f0 \'a0
\f1 \

\f0 \'a0
\f1 \

\f0 \'a0
\f1 \

\f0 \'a0
\f1 \

\f0 \'a0
\f1 \

\f0 \'a0
\f1 \

\f0 \'a0
\f1 \

\f0 \'a0
\f1 \

\f0 \'a0
\f1 \

\f0 \'a0
\f1 \

\f0 \'a0
\f1 \

\f0 \'a0
\f1 \

\f0 \'a0}